[aimspice]
[description]
921
excercie 4

*.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\�ving_4\p18_cmos_models_ss.inc
.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\�ving_4\p18_cmos_models_ff.inc
*.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\�ving_4\p18_cmos_models_tt.inc

.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\�ving_4\p18_model_card.inc

*MN1 DRAIN GATE SOURCE BULK WIDTH LENGTH
.subckt opampInverter Vin t

.param wn={0.9U}
.param L={0.18U}
.param wp={k*wn}
.param k=3.57

VDD vdd 0 dc 1.8v
*VIN Vin 0 dc 0.9v

MP1 t Vin vdd vdd PMOS L=0.18u W=wp
MN1 t Vin 0 0 NMOS L=0.18u W=wn

.ends 
xopamp1 1 2 opampInverter
xopamp2 2 3 opampInverter 
xopamp3 3 4 opampInverter 
xopamp4 4 5 opampInverter 
xopamp5 5 1 opampInverter

C1 1 0 100ff
C2 2 0 100ff
C3 3 0 100ff
C4 4 0 100ff
C5 5 0 100ff
.ic v(1)= 0.9v

.extract tran xdown(v(1,0.9<0100 ff,1000n>,100))
[tran]
0.1n
1000n
X
X
1
[ana]
4 1
0
1 1
1 1 0 5
1
v(1)
[end]

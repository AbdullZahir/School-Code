[aimspice]
[description]
1665
Analog circuit PROJECT(1 pixel)

.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\PROJECT\p18_cmos_models_tt.inc
.include C:\Users\Bruker\Documents\6_semester\Design_av_IC\PROJECT\p18_model_card.inc

*MN1 DRAIN GATE SOURCE BULK NMOS WIDTH LENGTH 
*MP1 SOURCE GATE DRAIN BULK PMOS WIDTH LENGTH
*0.7U<L<2U  2U<W<10U    Cs>=3pf    Cc1=Cc2=3pf   Vdd=1.8V

.param Wn={2u} 
.param Wp={2u}
.param Ln={0.7u}
.param Lp={0.7u}
.param Cs={3pf}
.param T=10

V_EXP gEXPOSE 0 PULSE(1.8 0 0 T/100 T/100 2 T)
V_ERASE gERASE  PULSE(0 1.8 0 T/100 T/100 2 T)

*gNRE (1.8 0 0 T/100 T/100 2 T) 
X1 
*-------------------------------------------------------------------------------------------------------------
.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 
*-------------------------------------------------------------------------------------------------------------
*F�rste delen av kretsen med nmos transistorer
.subckt  del_1 gEXPOSE gERASE vdd N1 N2 
*VDD-N1 
VDD1 vdd N1 dc 1.8v 
PhotoDiode vdd N1

*N1-N2
EXPOSE N1 gEXPOSE N2 0 NMOS L=Ln W=Wn
ERASE N2 gERASE 0 0 NMOS L=Ln W=Wn
CS N2 0 100ff
.ends 
*-------------------------------------------------------------------------------------------------------------
*Dette er andre delen av kretsen som best�r av pmos transistorer
.subckt del_2 N3 gNRE

MP3 N3 N2 0 vdd PMOS L=Lp W=Wp

*N3-OUT
NRE OUT gNRE N3 vdd PMOS L=Lp W=Wp
.ends
*-------------------------------------------------------------------------------------------------------------
x1 del_1


[tran]
0.1n
1000n
X
X
0
[ana]
4 0
[end]
